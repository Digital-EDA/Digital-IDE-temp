// Description: Package with constant APB v2.0 constants
package apb_pkg;

  typedef logic [2:0]  prot_t;

  localparam RESP_OKAY   = 1'b0;
  localparam RESP_SLVERR = 1'b1;

endpackage
